module InstructionMemory(Address, Instruction);
	input [31:0] Address;
	output reg [31:0] Instruction;
	
	always @(*)
		case (Address[9:2])
			8'd0: Instruction <= 32'h08000003;
			8'd1: Instruction <= 32'h08000067;
			8'd2: Instruction <= 32'h08000085;
			8'd3: Instruction <= 32'h201f0014;
			8'd4: Instruction <= 32'h03e00008;
			8'd5: Instruction <= 32'h3c174000;
			8'd6: Instruction <= 32'h8ef60014;
			8'd7: Instruction <= 32'h241d0400;
			8'd8: Instruction <= 32'h24040000;
			8'd9: Instruction <= 32'h24050000;
			8'd10: Instruction <= 32'h2406007f;
			8'd11: Instruction <= 32'h0c000022;
			8'd12: Instruction <= 32'h8ef50014;
			8'd13: Instruction <= 32'h02b6a022;
			8'd14: Instruction <= 32'h2408000f;
			8'd15: Instruction <= 32'h01148024;
			8'd16: Instruction <= 32'h0014a102;
			8'd17: Instruction <= 32'h01148824;
			8'd18: Instruction <= 32'h0014a102;
			8'd19: Instruction <= 32'h01149024;
			8'd20: Instruction <= 32'h0014a102;
			8'd21: Instruction <= 32'h01149824;
			8'd22: Instruction <= 32'h24080001;
			8'd23: Instruction <= 32'haee8000c;
			8'd24: Instruction <= 32'h24160000;
			8'd25: Instruction <= 32'h2001000f;
			8'd26: Instruction <= 32'h00014022;
			8'd27: Instruction <= 32'haee80000;
			8'd28: Instruction <= 32'h20010001;
			8'd29: Instruction <= 32'h00014022;
			8'd30: Instruction <= 32'haee80004;
			8'd31: Instruction <= 32'h24080003;
			8'd32: Instruction <= 32'haee80008;
			8'd33: Instruction <= 32'h08000021;
			8'd34: Instruction <= 32'h23bdfff0;
			8'd35: Instruction <= 32'hafbf000c;
			8'd36: Instruction <= 32'hafb20008;
			8'd37: Instruction <= 32'hafb10004;
			8'd38: Instruction <= 32'hafb00000;
			8'd39: Instruction <= 32'h00048021;
			8'd40: Instruction <= 32'h00058821;
			8'd41: Instruction <= 32'h00069021;
			8'd42: Instruction <= 32'h00114021;
			8'd43: Instruction <= 32'h00124821;
			8'd44: Instruction <= 32'h00115080;
			8'd45: Instruction <= 32'h020a5020;
			8'd46: Instruction <= 32'h8d530000;
			8'd47: Instruction <= 32'h00095080;
			8'd48: Instruction <= 32'h020a5020;
			8'd49: Instruction <= 32'h8d4b0000;
			8'd50: Instruction <= 32'h0173082b;
			8'd51: Instruction <= 32'h14200004;
			8'd52: Instruction <= 32'h0109082a;
			8'd53: Instruction <= 32'h10200002;
			8'd54: Instruction <= 32'h2129ffff;
			8'd55: Instruction <= 32'h0800002f;
			8'd56: Instruction <= 32'h00085080;
			8'd57: Instruction <= 32'h020a5020;
			8'd58: Instruction <= 32'h8d4b0000;
			8'd59: Instruction <= 32'h026b082b;
			8'd60: Instruction <= 32'h14200004;
			8'd61: Instruction <= 32'h0109082a;
			8'd62: Instruction <= 32'h10200002;
			8'd63: Instruction <= 32'h21080001;
			8'd64: Instruction <= 32'h08000038;
			8'd65: Instruction <= 32'h0109082a;
			8'd66: Instruction <= 32'h10200009;
			8'd67: Instruction <= 32'h00085080;
			8'd68: Instruction <= 32'h020a5020;
			8'd69: Instruction <= 32'h00095880;
			8'd70: Instruction <= 32'h020b5820;
			8'd71: Instruction <= 32'h8d4c0000;
			8'd72: Instruction <= 32'h8d6d0000;
			8'd73: Instruction <= 32'had6c0000;
			8'd74: Instruction <= 32'had4d0000;
			8'd75: Instruction <= 32'h0800002f;
			8'd76: Instruction <= 32'h00115080;
			8'd77: Instruction <= 32'h020a5020;
			8'd78: Instruction <= 32'h00085880;
			8'd79: Instruction <= 32'h020b5820;
			8'd80: Instruction <= 32'h8d6c0000;
			8'd81: Instruction <= 32'had4c0000;
			8'd82: Instruction <= 32'had730000;
			8'd83: Instruction <= 32'h210affff;
			8'd84: Instruction <= 32'h022a082a;
			8'd85: Instruction <= 32'h10200004;
			8'd86: Instruction <= 32'h00102021;
			8'd87: Instruction <= 32'h00112821;
			8'd88: Instruction <= 32'h000a3021;
			8'd89: Instruction <= 32'h0c000022;
			8'd90: Instruction <= 32'h210a0001;
			8'd91: Instruction <= 32'h0152082a;
			8'd92: Instruction <= 32'h10200004;
			8'd93: Instruction <= 32'h00102021;
			8'd94: Instruction <= 32'h000a2821;
			8'd95: Instruction <= 32'h00123021;
			8'd96: Instruction <= 32'h0c000022;
			8'd97: Instruction <= 32'h8fbf000c;
			8'd98: Instruction <= 32'h8fb20008;
			8'd99: Instruction <= 32'h8fb10004;
			8'd100: Instruction <= 32'h8fb00000;
			8'd101: Instruction <= 32'h23bd0010;
			8'd102: Instruction <= 32'h03e00008;
			8'd103: Instruction <= 32'h24080001;
			8'd104: Instruction <= 32'haee80008;
			8'd105: Instruction <= 32'h12c00009;
			8'd106: Instruction <= 32'h20010001;
			8'd107: Instruction <= 32'h02c14022;
			8'd108: Instruction <= 32'h11000009;
			8'd109: Instruction <= 32'h20010001;
			8'd110: Instruction <= 32'h01014022;
			8'd111: Instruction <= 32'h11000009;
			8'd112: Instruction <= 32'h20010001;
			8'd113: Instruction <= 32'h01014022;
			8'd114: Instruction <= 32'h11000009;
			8'd115: Instruction <= 32'h24080100;
			8'd116: Instruction <= 32'h01104020;
			8'd117: Instruction <= 32'h0800007f;
			8'd118: Instruction <= 32'h24080200;
			8'd119: Instruction <= 32'h01114020;
			8'd120: Instruction <= 32'h0800007f;
			8'd121: Instruction <= 32'h24080400;
			8'd122: Instruction <= 32'h01124020;
			8'd123: Instruction <= 32'h0800007f;
			8'd124: Instruction <= 32'h24080800;
			8'd125: Instruction <= 32'h01134020;
			8'd126: Instruction <= 32'h0800007f;
			8'd127: Instruction <= 32'h22d60001;
			8'd128: Instruction <= 32'h32d60003;
			8'd129: Instruction <= 32'haee80010;
			8'd130: Instruction <= 32'h24080003;
			8'd131: Instruction <= 32'haee80008;
			8'd132: Instruction <= 32'h03400008;
			8'd133: Instruction <= 32'h08000085;
			default: Instruction <= 32'h00000000;
		endcase
	
endmodule
